`timescale 1ns/1ns
module my_j1(input a0, b0, output j1);
	myXNOR G1(a0, b0, j1);
endmodule