`timescale 1ns/1ns
module threeB_counter_TB();
	logic clk = 0, en = 0;
	wire [2:0] po;
	wire co;
	threeB_counter TB1(clk, en, po, co);
	always #100 clk = ~clk;
	initial begin
	#150 en = ~en;
	#2000 $stop;
	end
endmodule